interface int_in;
  
  logic increment, reset, startstop, load;
  logic [1:0] digit_i;
  logic [3:0] value;
     
endinterface