package pkg_compilare;
  include "command.sv";
  include "generator.sv";
  include "driver.sv";
  include "monitor_input.sv";
  include "monitor_output.sv";
endpackage