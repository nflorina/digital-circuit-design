interface int_out;

  logic [6:0] cifra0, cifra1, cifra2, cifra3;
     
endinterface